module basic_module (input clk,
input rst,
output [7:0] data);
wire [15:0] internal_signal;
reg [31:0] counter;
endmodule